* C:\Users\Lenovo\eSim-Workspace\test\test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 02/01/25 10:46:42

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  out in GND GND mosfet_n		
M2  Net-_M2-Pad1_ in out Net-_M2-Pad1_ mosfet_p		
v2  Net-_M2-Pad1_ GND DC		
v1  in GND pulse		
U1  in plot_v1		
U2  out plot_v1		

.end
