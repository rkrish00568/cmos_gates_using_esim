* C:\Users\Lenovo\eSim-Workspace\nanddd\nanddd.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 02/08/25 20:05:25

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M2  Vout Ain Net-_M2-Pad3_ GND eSim_MOS_N		
M1  Net-_M1-Pad1_ Ain Vout Net-_M1-Pad1_ eSim_MOS_P		
v3  Net-_M1-Pad1_ GND DC		
M3  Net-_M2-Pad3_ Bin GND GND eSim_MOS_N		
v2  Bin GND pulse		
v1  Ain GND pulse		
M4  Net-_M1-Pad1_ Bin Vout Net-_M1-Pad1_ eSim_MOS_P		
U1  Ain plot_v1		
U2  Bin plot_v1		
U3  Vout plot_v1		

.end
