* C:\Users\Lenovo\eSim-Workspace\or_with_nansd\or_with_nansd.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 02/27/25 11:26:05

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U2-Pad1_ Net-_U2-Pad1_ Net-_U2-Pad3_ d_nand		
v1  in GND pulse		
U3  out plot_v1		
U1  in plot_v1		
U4  in Net-_U2-Pad1_ adc_bridge_1		
U5  Net-_U2-Pad3_ out dac_bridge_1		

.end
